module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_Counter # (.UUID(64'd2452350458780268905 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_0 (.clk(clk), .rst(rst), .save(wire_98), .in(wire_0), .out(wire_102));
  TC_Splitter8 # (.UUID(64'd1580408133110145864 ^ UUID)) Splitter8_1 (.in(wire_46[7:0]), .out0(wire_57), .out1(wire_120), .out2(wire_68), .out3(), .out4(wire_75), .out5(wire_78), .out6(wire_65), .out7(wire_81));
  TC_Splitter8 # (.UUID(64'd2059178242977121373 ^ UUID)) Splitter8_2 (.in(wire_12[7:0]), .out0(wire_114), .out1(wire_113), .out2(wire_116), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2693264835291803615 ^ UUID)) Splitter8_3 (.in(wire_101[7:0]), .out0(wire_122), .out1(wire_109), .out2(wire_60), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd158812426551174434 ^ UUID)) Splitter8_4 (.in(wire_77[7:0]), .out0(wire_79), .out1(wire_42), .out2(wire_40), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3092528147277599578 ^ UUID)) Decoder3_5 (.dis(wire_41), .sel0(wire_79), .sel1(wire_42), .sel2(wire_40), .out0(wire_73), .out1(wire_100), .out2(wire_58), .out3(wire_104), .out4(wire_96), .out5(wire_13), .out6(wire_83), .out7(wire_124));
  TC_Decoder3 # (.UUID(64'd2474399514938988928 ^ UUID)) Decoder3_6 (.dis(wire_81), .sel0(wire_114), .sel1(wire_113), .sel2(wire_116), .out0(wire_7), .out1(wire_36), .out2(wire_32), .out3(wire_85), .out4(wire_43), .out5(wire_92), .out6(), .out7(wire_33));
  TC_Decoder3 # (.UUID(64'd806511425691535975 ^ UUID)) Decoder3_7 (.dis(wire_65), .sel0(wire_122), .sel1(wire_109), .sel2(wire_60), .out0(wire_70), .out1(wire_1), .out2(wire_9), .out3(wire_55), .out4(wire_8), .out5(wire_10), .out6(), .out7(wire_5));
  TC_IOSwitch # (.UUID(64'd4186197826621441477 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_8 (.in(wire_11), .en(wire_124), .out(arch_output_value));
  TC_Switch # (.UUID(64'd3276341372597245191 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_9 (.en(wire_54), .in(arch_input_value), .out(wire_31));
  TC_Or # (.UUID(64'd2926217265011126760 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_7), .in1(wire_70), .out(wire_59));
  TC_Or # (.UUID(64'd4346183087953155811 ^ UUID), .BIT_WIDTH(64'd1)) Or_11 (.in0(wire_36), .in1(wire_1), .out(wire_103));
  TC_Or # (.UUID(64'd134634696612420425 ^ UUID), .BIT_WIDTH(64'd1)) Or_12 (.in0(wire_32), .in1(wire_9), .out(wire_27));
  TC_Or # (.UUID(64'd1969669177385825140 ^ UUID), .BIT_WIDTH(64'd1)) Or_13 (.in0(wire_85), .in1(wire_55), .out(wire_90));
  TC_Or # (.UUID(64'd2125493594201118714 ^ UUID), .BIT_WIDTH(64'd1)) Or_14 (.in0(wire_43), .in1(wire_8), .out(wire_35));
  TC_Switch # (.UUID(64'd3578892536211673484 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_7), .in(wire_107), .out(wire_16_0));
  TC_Switch # (.UUID(64'd1560654892581336712 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_36), .in(wire_19), .out(wire_16_1));
  TC_Switch # (.UUID(64'd1811287876483295164 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_32), .in(wire_66), .out(wire_16_2));
  TC_Switch # (.UUID(64'd2080533949957218959 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_70), .in(wire_107), .out(wire_24_6));
  TC_Switch # (.UUID(64'd3382407185197042630 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_1), .in(wire_19), .out(wire_24_5));
  TC_Switch # (.UUID(64'd1899559205710328747 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_5), .in(wire_31), .out(wire_24_0));
  TC_Switch # (.UUID(64'd4577499525846200431 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_33), .in(wire_31), .out(wire_16_6));
  TC_Switch # (.UUID(64'd2151517462767163191 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_9), .in(wire_66), .out(wire_24_4));
  TC_Switch # (.UUID(64'd4194123250794237968 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_85), .in(wire_126), .out(wire_16_3));
  TC_Switch # (.UUID(64'd1353324206004192233 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_55), .in(wire_126), .out(wire_24_3));
  TC_Switch # (.UUID(64'd844909057701417619 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_43), .in(wire_25), .out(wire_16_5));
  TC_Switch # (.UUID(64'd3267461772374150223 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_8), .in(wire_25), .out(wire_24_2));
  TC_Or # (.UUID(64'd753993920865946244 ^ UUID), .BIT_WIDTH(64'd1)) Or_27 (.in0(wire_33), .in1(wire_5), .out(wire_54));
  TC_Register # (.UUID(64'd1473628890728886837 ^ UUID), .BIT_WIDTH(64'd8)) Register8_28 (.clk(clk), .rst(rst), .load(wire_59), .save(wire_73), .in(wire_11), .out(wire_107));
  TC_Register # (.UUID(64'd3404127598317107480 ^ UUID), .BIT_WIDTH(64'd8)) Register8_29 (.clk(clk), .rst(rst), .load(wire_103), .save(wire_100), .in(wire_11), .out(wire_19));
  TC_Register # (.UUID(64'd857710086233477403 ^ UUID), .BIT_WIDTH(64'd8)) Register8_30 (.clk(clk), .rst(rst), .load(wire_27), .save(wire_58), .in(wire_11), .out(wire_66));
  TC_Register # (.UUID(64'd716496557207202822 ^ UUID), .BIT_WIDTH(64'd8)) Register8_31 (.clk(clk), .rst(rst), .load(wire_90), .save(wire_104), .in(wire_11), .out(wire_126));
  TC_Register # (.UUID(64'd4308546724317967359 ^ UUID), .BIT_WIDTH(64'd8)) Register8_32 (.clk(clk), .rst(rst), .load(wire_35), .save(wire_96), .in(wire_11), .out(wire_25));
  TC_Or # (.UUID(64'd1131191003299457672 ^ UUID), .BIT_WIDTH(64'd8)) Or8_33 (.in0(wire_106), .in1(wire_24), .out(wire_2));
  TC_Or # (.UUID(64'd3658741303214134569 ^ UUID), .BIT_WIDTH(64'd8)) Or8_34 (.in0(wire_94), .in1(wire_16), .out(wire_4));
  TC_Switch # (.UUID(64'd2531986671109172071 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_65), .in(wire_101[7:0]), .out(wire_106));
  TC_Switch # (.UUID(64'd829754361863765621 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_36 (.en(wire_81), .in(wire_12[7:0]), .out(wire_94));
  TC_Switch # (.UUID(64'd3809920487273635419 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_37 (.en(wire_92), .in(wire_18), .out(wire_16_4));
  TC_Switch # (.UUID(64'd4089127036144108990 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_38 (.en(wire_10), .in(wire_18), .out(wire_24_1));
  TC_Or # (.UUID(64'd3539695120833480884 ^ UUID), .BIT_WIDTH(64'd1)) Or_39 (.in0(wire_92), .in1(wire_10), .out(wire_63));
  TC_Decoder3 # (.UUID(64'd959215858486299202 ^ UUID)) Decoder3_40 (.dis(1'd0), .sel0(wire_57), .sel1(wire_120), .sel2(wire_68), .out0(wire_119), .out1(wire_111), .out2(wire_39), .out3(wire_110), .out4(wire_112), .out5(wire_62), .out6(wire_131), .out7(wire_125));
  TC_Add # (.UUID(64'd488376956936131461 ^ UUID), .BIT_WIDTH(64'd8)) Add8_41 (.in0(wire_4), .in1(wire_2), .ci(1'd0), .out(wire_95), .co());
  TC_Switch # (.UUID(64'd4121249633311310994 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_42 (.en(wire_72), .in(wire_95), .out(wire_3_2));
  TC_Neg # (.UUID(64'd4540844933532444684 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_43 (.in(wire_2), .out(wire_76));
  TC_Add # (.UUID(64'd945362313428989074 ^ UUID), .BIT_WIDTH(64'd8)) Add8_44 (.in0(wire_4), .in1(wire_76), .ci(1'd0), .out(wire_118), .co());
  TC_Switch # (.UUID(64'd1130487566684413615 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_44), .in(wire_118), .out(wire_3_0));
  TC_Maker8 # (.UUID(64'd3552730175243824440 ^ UUID)) Maker8_46 (.in0(wire_119), .in1(wire_111), .in2(wire_39), .in3(wire_110), .in4(wire_112), .in5(wire_62), .in6(wire_131), .in7(wire_125), .out(wire_61));
  TC_Splitter8 # (.UUID(64'd462425196375030397 ^ UUID)) Splitter8_47 (.in(wire_61), .out0(wire_72), .out1(wire_44), .out2(wire_48), .out3(wire_56), .out4(wire_91), .out5(wire_64), .out6(wire_105), .out7(wire_97));
  TC_Switch # (.UUID(64'd2403089770491926697 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_74), .in(wire_3), .out(wire_11_0));
  TC_And # (.UUID(64'd2149687390567888029 ^ UUID), .BIT_WIDTH(64'd8)) And8_49 (.in0(wire_4), .in1(wire_2), .out(wire_67));
  TC_Or # (.UUID(64'd3471921671444333826 ^ UUID), .BIT_WIDTH(64'd8)) Or8_50 (.in0(wire_4), .in1(wire_2), .out(wire_99));
  TC_Not # (.UUID(64'd689544037905960133 ^ UUID), .BIT_WIDTH(64'd8)) Not8_51 (.in(wire_4), .out(wire_123));
  TC_Xor # (.UUID(64'd2961167983726257251 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_52 (.in0(wire_4), .in1(wire_2), .out(wire_52));
  TC_Switch # (.UUID(64'd4559915573104512857 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_48), .in(wire_67), .out(wire_3_1));
  TC_Switch # (.UUID(64'd90038848783738937 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_56), .in(wire_99), .out(wire_3_3));
  TC_Switch # (.UUID(64'd2551781636376953774 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_55 (.en(wire_91), .in(wire_123), .out(wire_3_4));
  TC_Switch # (.UUID(64'd2046784265305930612 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_56 (.en(wire_64), .in(wire_52), .out(wire_3_5));
  TC_Mul # (.UUID(64'd2211514518710572405 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_57 (.in0(wire_4), .in1(wire_2), .out0(wire_30), .out1(wire_127));
  TC_Switch # (.UUID(64'd198050465957076576 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_58 (.en(wire_97), .in(wire_127), .out(wire_3_7));
  TC_Switch # (.UUID(64'd2712460921153961372 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_59 (.en(wire_105), .in(wire_30), .out(wire_3_6));
  TC_Splitter8 # (.UUID(64'd951832874730727267 ^ UUID)) Splitter8_60 (.in(wire_61), .out0(wire_88), .out1(wire_29), .out2(wire_20), .out3(wire_86), .out4(wire_37), .out5(wire_71), .out6(wire_108), .out7(wire_17));
  TC_Equal # (.UUID(64'd2298929716682680619 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_61 (.in0(wire_4), .in1(wire_2), .out(wire_47));
  TC_Switch # (.UUID(64'd4182284540579803752 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_62 (.en(wire_88), .in(wire_47), .out(wire_14_4));
  TC_Not # (.UUID(64'd662622555333555876 ^ UUID), .BIT_WIDTH(64'd1)) Not_63 (.in(wire_47), .out(wire_93));
  TC_Switch # (.UUID(64'd1438853858099742271 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_64 (.en(wire_29), .in(wire_93), .out(wire_14_2));
  TC_LessU # (.UUID(64'd523447668447656097 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_65 (.in0(wire_4), .in1(wire_2), .out(wire_22));
  TC_Switch # (.UUID(64'd2407577354869023759 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_66 (.en(wire_20), .in(wire_22), .out(wire_14_0));
  TC_Or # (.UUID(64'd865387050054296889 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_22), .in1(wire_47), .out(wire_132));
  TC_Switch # (.UUID(64'd3430743913552632765 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_68 (.en(wire_86), .in(wire_132), .out(wire_14_1));
  TC_Nor # (.UUID(64'd4472183732922582580 ^ UUID), .BIT_WIDTH(64'd1)) Nor_69 (.in0(wire_22), .in1(wire_47), .out(wire_129));
  TC_Switch # (.UUID(64'd3306992519549871553 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_70 (.en(wire_37), .in(wire_129), .out(wire_14_3));
  TC_Not # (.UUID(64'd2955059209242120201 ^ UUID), .BIT_WIDTH(64'd1)) Not_71 (.in(wire_22), .out(wire_26));
  TC_Switch # (.UUID(64'd3227335121701824192 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_72 (.en(wire_71), .in(wire_26), .out(wire_14_5));
  TC_Switch # (.UUID(64'd2683517932211923067 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_73 (.en(wire_15), .in(wire_14), .out(wire_41));
  TC_Mul # (.UUID(64'd2563314739157226883 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_74 (.in0(wire_4), .in1(wire_45), .out0(wire_121), .out1(wire_89));
  TC_Switch # (.UUID(64'd3929656369738992149 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_108), .in(wire_121), .out(wire_6_0));
  TC_Switch # (.UUID(64'd3063638702614327857 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_76 (.en(wire_17), .in(wire_89), .out(wire_6_1));
  TC_Switch # (.UUID(64'd4553200895106409104 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_77 (.en(wire_15), .in(wire_6), .out(wire_11_1));
  TC_Mux # (.UUID(64'd791295078858124393 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_78 (.sel(wire_115), .in0({{7{1'b0}}, wire_128 }), .in1(wire_2), .out(wire_45));
  TC_Constant # (.UUID(64'd4510222432388480606 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_79 (.out(wire_128));
  TC_Or # (.UUID(64'd1015712669360850097 ^ UUID), .BIT_WIDTH(64'd1)) Or_80 (.in0(wire_108), .in1(wire_17), .out(wire_115));
  TC_Mux # (.UUID(64'd2625454164047475578 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_81 (.sel(wire_41), .in0(wire_11), .in1(wire_77[7:0]), .out(wire_0));
  TC_Or # (.UUID(64'd2168341804967303507 ^ UUID), .BIT_WIDTH(64'd1)) Or_82 (.in0(wire_83), .in1(wire_41), .out(wire_98));
  TC_Splitter8 # (.UUID(64'd1290519562063653211 ^ UUID)) Splitter8_83 (.in(wire_61), .out0(wire_87), .out1(wire_82), .out2(wire_80), .out3(wire_51), .out4(wire_38), .out5(wire_50), .out6(wire_53), .out7());
  TC_Ashr # (.UUID(64'd846670947147293708 ^ UUID), .BIT_WIDTH(64'd8)) Ashr8_84 (.in(wire_4), .shift(wire_2), .out(wire_69));
  TC_Ror # (.UUID(64'd2902599177739172371 ^ UUID), .BIT_WIDTH(64'd8)) Ror8_85 (.in(wire_4), .shift(wire_2), .out(wire_49));
  TC_Rol # (.UUID(64'd3040107488757936910 ^ UUID), .BIT_WIDTH(64'd8)) Rol8_86 (.in(wire_4), .shift(wire_2), .out(wire_34));
  TC_Shr # (.UUID(64'd3261478892196693155 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_87 (.in(wire_4), .shift(wire_2), .out(wire_117));
  TC_Shl # (.UUID(64'd3163731994518766222 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_88 (.in(wire_4), .shift(wire_2), .out(wire_130));
  TC_Switch # (.UUID(64'd587093708640519058 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_89 (.en(wire_87), .in(wire_69), .out(wire_21_0));
  TC_Switch # (.UUID(64'd218368253074601695 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_90 (.en(wire_82), .in(wire_49), .out(wire_21_1));
  TC_Switch # (.UUID(64'd1164417289337729766 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_91 (.en(wire_80), .in(wire_34), .out(wire_21_2));
  TC_Switch # (.UUID(64'd339117104162153763 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_92 (.en(wire_51), .in(wire_117), .out(wire_21_3));
  TC_Switch # (.UUID(64'd345196551137786680 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_93 (.en(wire_38), .in(wire_130), .out(wire_21_4));
  TC_Switch # (.UUID(64'd1967651675007569350 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_94 (.en(wire_23), .in(wire_21), .out(wire_11_2));
  TC_Ram # (.UUID(64'd773551801835591906 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_95 (.clk(clk), .rst(rst), .load(wire_50), .save(wire_53), .address({{24{1'b0}}, wire_28 }), .in0({{56{1'b0}}, wire_4 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_84), .out1(), .out2(), .out3());
  TC_Switch # (.UUID(64'd200221941951721592 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_96 (.en(wire_50), .in(wire_84[7:0]), .out(wire_11_3));
  _2z_bitz_decoder # (.UUID(64'd4345311738281130334 ^ UUID)) _2z_bitz_decoder_97 (.clk(clk), .rst(rst), .Input_1(wire_75), .Input_2(wire_78), .Output_1(wire_74), .Output_2(), .Output_3(wire_23), .Output_4(wire_15));
  RegisterPlus # (.UUID(64'd336705455147415054 ^ UUID)) RegisterPlus_98 (.clk(clk), .rst(rst), .Load(wire_63), .Save_value(wire_11), .Save(wire_13), .Always_output(wire_28), .Output(wire_18));
  TC_Program # (.UUID(64'd1403467390952442459 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_137A1E27FB908A5B.w8.bin"), .ARG_SIG("Program_137A1E27FB908A5B=%s")) Program_99 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_102 }), .out0(wire_46), .out1(wire_12), .out2(wire_101), .out3(wire_77));

  wire [7:0] wire_0;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  wire [7:0] wire_3_2;
  wire [7:0] wire_3_3;
  wire [7:0] wire_3_4;
  wire [7:0] wire_3_5;
  wire [7:0] wire_3_6;
  wire [7:0] wire_3_7;
  assign wire_3 = wire_3_0|wire_3_1|wire_3_2|wire_3_3|wire_3_4|wire_3_5|wire_3_6|wire_3_7;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_6_0;
  wire [7:0] wire_6_1;
  assign wire_6 = wire_6_0|wire_6_1;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_11_0;
  wire [7:0] wire_11_1;
  wire [7:0] wire_11_2;
  wire [7:0] wire_11_3;
  assign wire_11 = wire_11_0|wire_11_1|wire_11_2|wire_11_3;
  wire [63:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_14_0;
  wire [0:0] wire_14_1;
  wire [0:0] wire_14_2;
  wire [0:0] wire_14_3;
  wire [0:0] wire_14_4;
  wire [0:0] wire_14_5;
  assign wire_14 = wire_14_0|wire_14_1|wire_14_2|wire_14_3|wire_14_4|wire_14_5;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_16_0;
  wire [7:0] wire_16_1;
  wire [7:0] wire_16_2;
  wire [7:0] wire_16_3;
  wire [7:0] wire_16_4;
  wire [7:0] wire_16_5;
  wire [7:0] wire_16_6;
  assign wire_16 = wire_16_0|wire_16_1|wire_16_2|wire_16_3|wire_16_4|wire_16_5|wire_16_6;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [7:0] wire_21_0;
  wire [7:0] wire_21_1;
  wire [7:0] wire_21_2;
  wire [7:0] wire_21_3;
  wire [7:0] wire_21_4;
  assign wire_21 = wire_21_0|wire_21_1|wire_21_2|wire_21_3|wire_21_4;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_24_0;
  wire [7:0] wire_24_1;
  wire [7:0] wire_24_2;
  wire [7:0] wire_24_3;
  wire [7:0] wire_24_4;
  wire [7:0] wire_24_5;
  wire [7:0] wire_24_6;
  assign wire_24 = wire_24_0|wire_24_1|wire_24_2|wire_24_3|wire_24_4|wire_24_5|wire_24_6;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [7:0] wire_45;
  wire [63:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [7:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  assign arch_input_enable = wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [7:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [7:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [7:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [7:0] wire_76;
  wire [63:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [63:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [7:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [7:0] wire_94;
  wire [7:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [7:0] wire_99;
  wire [0:0] wire_100;
  wire [63:0] wire_101;
  wire [7:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [7:0] wire_106;
  wire [7:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [7:0] wire_117;
  wire [7:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [7:0] wire_121;
  wire [0:0] wire_122;
  wire [7:0] wire_123;
  wire [0:0] wire_124;
  assign arch_output_enable = wire_124;
  wire [0:0] wire_125;
  wire [7:0] wire_126;
  wire [7:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [7:0] wire_130;
  wire [0:0] wire_131;
  wire [0:0] wire_132;

endmodule
